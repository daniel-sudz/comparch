`timescale 1ns/1ps
`default_nettype none


/* Sample file to compile */

module sample (input logic a, output logic b);
    assign b = a;
endmodule