/*
 * Header Information
 *
 */

module simple_in_n_out (in_1,
                        in_2,
                        in_3);
    
    /* Port definition */
    input in_1;
    input in_2;
    input in_3;
    
    
endmodule
